//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Fri Jun 04 10:12:51 2021
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// TPLSRAM_32x512BIT
module TPLSRAM_32x512BIT(
    // Inputs
    RADDR,
    RCLK,
    WADDR,
    WCLK,
    WD,
    WEN,
    // Outputs
    RD
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  [8:0]  RADDR;
input         RCLK;
input  [8:0]  WADDR;
input         WCLK;
input  [31:0] WD;
input         WEN;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [31:0] RD;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   [8:0]  RADDR;
wire          RCLK;
wire   [31:0] RD_0;
wire   [8:0]  WADDR;
wire          WCLK;
wire   [31:0] WD;
wire          WEN;
wire   [31:0] RD_0_net_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire          GND_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net = 1'b0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign RD_0_net_0 = RD_0;
assign RD[31:0]   = RD_0_net_0;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------TPLSRAM_32x512BIT_TPLSRAM_32x512BIT_0_TPSRAM   -   Actel:SgCore:TPSRAM:1.0.101
TPLSRAM_32x512BIT_TPLSRAM_32x512BIT_0_TPSRAM TPLSRAM_32x512BIT_0(
        // Inputs
        .WEN   ( WEN ),
        .WCLK  ( WCLK ),
        .RCLK  ( RCLK ),
        .WD    ( WD ),
        .WADDR ( WADDR ),
        .RADDR ( RADDR ),
        // Outputs
        .RD    ( RD_0 ) 
        );


endmodule
