library verilog;
use verilog.vl_types.all;
entity AHBLite_CAN_Bridge is
    generic(
        AHB_Lite_FSM_Get_ADDR: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Get_Data_2_CAN_A: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        AHB_Lite_FSM_Get_Data_2_CAN_B: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        AHB_Lite_FSM_Get_Data_2_CAN_C: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        AHB_Lite_FSM_Get_Data_2_CAN_D: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Wait_CAN_A_Write: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Wait_CAN_B_Write: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Wait_CAN_C_Write: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Wait_CAN_D_Write: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Wait_CAN_A_Read: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Wait_CAN_B_Read: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Wait_CAN_C_Read: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Wait_CAN_D_Read: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Send_Data: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Read_Addr_Err: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        HREADYOUT_RDY   : vl_logic := Hi1;
        HREADYOUT_BSY   : vl_logic := Hi0;
        HRESP_OKAY      : vl_logic := Hi0;
        CAN_Operate_FSM_IDLE: integer := 0;
        CAN_Operate_FSM_A_Latch_ADDR_1st: integer := 1;
        CAN_Operate_FSM_A_Latch_ADDR_2nd: integer := 2;
        CAN_Operate_FSM_A_Read_Data_1st: integer := 4;
        CAN_Operate_FSM_A_Read_Data_2nd: integer := 8;
        CAN_Operate_FSM_A_Read_Data_3rd: integer := 16;
        CAN_Operate_FSM_A_Write_Data_1st: integer := 32;
        CAN_Operate_FSM_A_Write_Data_2nd: integer := 64;
        CAN_Operate_FSM_B_Latch_ADDR_1st: integer := 128;
        CAN_Operate_FSM_B_Latch_ADDR_2nd: integer := 256;
        CAN_Operate_FSM_B_Read_Data_1st: integer := 512;
        CAN_Operate_FSM_B_Read_Data_2nd: integer := 1024;
        CAN_Operate_FSM_B_Read_Data_3rd: integer := 2048;
        CAN_Operate_FSM_B_Write_Data_1st: integer := 4096;
        CAN_Operate_FSM_B_Write_Data_2nd: integer := 8192;
        CAN_Operate_FSM_C_Latch_ADDR_1st: integer := 16384;
        CAN_Operate_FSM_C_Latch_ADDR_2nd: integer := 32768;
        CAN_Operate_FSM_C_Read_Data_1st: integer := 65536;
        CAN_Operate_FSM_C_Read_Data_2nd: integer := 131072;
        CAN_Operate_FSM_C_Read_Data_3rd: integer := 262144;
        CAN_Operate_FSM_C_Write_Data_1st: integer := 524288;
        CAN_Operate_FSM_C_Write_Data_2nd: integer := 1048576;
        CAN_Operate_FSM_D_Latch_ADDR_1st: integer := 2097152;
        CAN_Operate_FSM_D_Latch_ADDR_2nd: integer := 4194304;
        CAN_Operate_FSM_D_Read_Data_1st: integer := 8388608;
        CAN_Operate_FSM_D_Read_Data_2nd: integer := 16777216;
        CAN_Operate_FSM_D_Read_Data_3rd: integer := 33554432;
        CAN_Operate_FSM_D_Write_Data_1st: integer := 67108864;
        CAN_Operate_FSM_D_Write_Data_2nd: integer := 134217728;
        CAN_Operate_FSM_Over: integer := 268435456;
        CAN_PORT_DIR_OUT: vl_logic := Hi0;
        CAN_PORT_DIR_IN : vl_logic := Hi1
    );
    port(
        HRESETn         : in     vl_logic;
        HCLK            : in     vl_logic;
        HSEL            : in     vl_logic;
        HADDR           : in     vl_logic_vector(31 downto 0);
        HWRITE          : in     vl_logic;
        HSIZE           : in     vl_logic_vector(2 downto 0);
        HBURST          : in     vl_logic_vector(2 downto 0);
        HPROT           : in     vl_logic_vector(3 downto 0);
        HTRANS          : in     vl_logic_vector(1 downto 0);
        HMASTLOCK       : in     vl_logic;
        HREADY          : in     vl_logic;
        HWDATA          : in     vl_logic_vector(31 downto 0);
        HRDATA          : out    vl_logic_vector(31 downto 0);
        HREADYOUT       : out    vl_logic;
        HRESP           : out    vl_logic;
        CAN_CLK         : in     vl_logic;
        CAN_RST         : out    vl_logic;
        CAN_A_ALE       : out    vl_logic;
        CAN_A_RD        : out    vl_logic;
        CAN_A_WR        : out    vl_logic;
        CAN_A_CS        : out    vl_logic;
        CAN_A_Port      : inout  vl_logic_vector(7 downto 0);
        CAN_B_ALE       : out    vl_logic;
        CAN_B_RD        : out    vl_logic;
        CAN_B_WR        : out    vl_logic;
        CAN_B_CS        : out    vl_logic;
        CAN_B_Port      : inout  vl_logic_vector(7 downto 0);
        CAN_C_ALE       : out    vl_logic;
        CAN_C_RD        : out    vl_logic;
        CAN_C_WR        : out    vl_logic;
        CAN_C_CS        : out    vl_logic;
        CAN_C_Port      : inout  vl_logic_vector(7 downto 0);
        CAN_D_ALE       : out    vl_logic;
        CAN_D_RD        : out    vl_logic;
        CAN_D_WR        : out    vl_logic;
        CAN_D_CS        : out    vl_logic;
        CAN_D_Port      : inout  vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Get_ADDR : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Get_Data_2_CAN_A : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Get_Data_2_CAN_B : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Get_Data_2_CAN_C : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Get_Data_2_CAN_D : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Wait_CAN_A_Write : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Wait_CAN_B_Write : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Wait_CAN_C_Write : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Wait_CAN_D_Write : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Wait_CAN_A_Read : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Wait_CAN_B_Read : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Wait_CAN_C_Read : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Wait_CAN_D_Read : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Send_Data : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Read_Addr_Err : constant is 1;
    attribute mti_svvh_generic_type of HREADYOUT_RDY : constant is 1;
    attribute mti_svvh_generic_type of HREADYOUT_BSY : constant is 1;
    attribute mti_svvh_generic_type of HRESP_OKAY : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_IDLE : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_A_Latch_ADDR_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_A_Latch_ADDR_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_A_Read_Data_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_A_Read_Data_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_A_Read_Data_3rd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_A_Write_Data_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_A_Write_Data_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_B_Latch_ADDR_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_B_Latch_ADDR_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_B_Read_Data_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_B_Read_Data_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_B_Read_Data_3rd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_B_Write_Data_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_B_Write_Data_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_C_Latch_ADDR_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_C_Latch_ADDR_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_C_Read_Data_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_C_Read_Data_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_C_Read_Data_3rd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_C_Write_Data_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_C_Write_Data_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_D_Latch_ADDR_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_D_Latch_ADDR_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_D_Read_Data_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_D_Read_Data_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_D_Read_Data_3rd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_D_Write_Data_1st : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_D_Write_Data_2nd : constant is 1;
    attribute mti_svvh_generic_type of CAN_Operate_FSM_Over : constant is 1;
    attribute mti_svvh_generic_type of CAN_PORT_DIR_OUT : constant is 1;
    attribute mti_svvh_generic_type of CAN_PORT_DIR_IN : constant is 1;
end AHBLite_CAN_Bridge;
