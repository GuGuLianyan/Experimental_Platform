library verilog;
use verilog.vl_types.all;
entity CLKINT_PRESERVE is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end CLKINT_PRESERVE;
