library verilog;
use verilog.vl_types.all;
entity bridge_tb is
end bridge_tb;
