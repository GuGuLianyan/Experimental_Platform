library verilog;
use verilog.vl_types.all;
entity AHBLite_1553_Bridge is
    generic(
        Interrupt_Mask_reg_RW: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        Config_reg_1_RW : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        Config_reg_2_RW : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        Start_Reset_reg_WO: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        RT_CMD_Stack_Point_reg_RO: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        RT_SubAddr_CTRL_Word_reg_RW: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        TimeScale_reg_RW: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        Interrupt_State_reg_RO: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        Config_reg_3_RW : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        Config_reg_4_RW : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        Config_reg_5_RW : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        RT_Data_Stack_Addr_reg_RW: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        RT_Last_CMD_Word_reg_RW: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        RT_State_Word_reg_RO: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        RT_BIT_reg_RO   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        AHB_Lite_FSM_Get_ADDR: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AHB_Lite_FSM_Get_Data: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        AHB_Lite_FSM_Wait_1553_Write: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        AHB_Lite_FSM_Wait_1553_Read: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        AHB_Lite_FSM_Send_Data: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        HREADYOUT_RDY   : vl_logic := Hi1;
        HREADYOUT_BSY   : vl_logic := Hi0;
        HRESP_OKAY      : vl_logic := Hi0;
        B1553_FSM_IDLE  : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        B1553_FSM_CS    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        B1553_FSM_Write : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        B1553_FSM_Read  : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        B1553_FSM_Wait_RDY: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        B1553_FSM_Over  : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        B1553_DATA_DIR_IN: vl_logic := Hi0;
        B1553_DATA_DIR_OUT: vl_logic := Hi1
    );
    port(
        HRESETn         : in     vl_logic;
        HCLK            : in     vl_logic;
        HSEL            : in     vl_logic;
        HADDR           : in     vl_logic_vector(31 downto 0);
        HWRITE          : in     vl_logic;
        HSIZE           : in     vl_logic_vector(2 downto 0);
        HBURST          : in     vl_logic_vector(2 downto 0);
        HPROT           : in     vl_logic_vector(3 downto 0);
        HTRANS          : in     vl_logic_vector(1 downto 0);
        HMASTLOCK       : in     vl_logic;
        HREADY          : in     vl_logic;
        HWDATA          : in     vl_logic_vector(31 downto 0);
        HRDATA          : out    vl_logic_vector(31 downto 0);
        HREADYOUT       : out    vl_logic;
        HRESP           : out    vl_logic;
        B1553_DATA_DIR  : out    vl_logic;
        CLK_16MHz       : in     vl_logic;
        B1553_ADDR      : out    vl_logic_vector(11 downto 0);
        B1553_DATA      : inout  vl_logic_vector(15 downto 0);
        B1553_RSTn      : out    vl_logic;
        B1553_CSn       : out    vl_logic;
        B1553_MEM_REGn  : out    vl_logic;
        B1553_RD_WRn    : out    vl_logic;
        B1553_RDYn      : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of Interrupt_Mask_reg_RW : constant is 1;
    attribute mti_svvh_generic_type of Config_reg_1_RW : constant is 1;
    attribute mti_svvh_generic_type of Config_reg_2_RW : constant is 1;
    attribute mti_svvh_generic_type of Start_Reset_reg_WO : constant is 1;
    attribute mti_svvh_generic_type of RT_CMD_Stack_Point_reg_RO : constant is 1;
    attribute mti_svvh_generic_type of RT_SubAddr_CTRL_Word_reg_RW : constant is 1;
    attribute mti_svvh_generic_type of TimeScale_reg_RW : constant is 1;
    attribute mti_svvh_generic_type of Interrupt_State_reg_RO : constant is 1;
    attribute mti_svvh_generic_type of Config_reg_3_RW : constant is 1;
    attribute mti_svvh_generic_type of Config_reg_4_RW : constant is 1;
    attribute mti_svvh_generic_type of Config_reg_5_RW : constant is 1;
    attribute mti_svvh_generic_type of RT_Data_Stack_Addr_reg_RW : constant is 1;
    attribute mti_svvh_generic_type of RT_Last_CMD_Word_reg_RW : constant is 1;
    attribute mti_svvh_generic_type of RT_State_Word_reg_RO : constant is 1;
    attribute mti_svvh_generic_type of RT_BIT_reg_RO : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Get_ADDR : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Get_Data : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Wait_1553_Write : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Wait_1553_Read : constant is 1;
    attribute mti_svvh_generic_type of AHB_Lite_FSM_Send_Data : constant is 1;
    attribute mti_svvh_generic_type of HREADYOUT_RDY : constant is 1;
    attribute mti_svvh_generic_type of HREADYOUT_BSY : constant is 1;
    attribute mti_svvh_generic_type of HRESP_OKAY : constant is 1;
    attribute mti_svvh_generic_type of B1553_FSM_IDLE : constant is 1;
    attribute mti_svvh_generic_type of B1553_FSM_CS : constant is 1;
    attribute mti_svvh_generic_type of B1553_FSM_Write : constant is 1;
    attribute mti_svvh_generic_type of B1553_FSM_Read : constant is 1;
    attribute mti_svvh_generic_type of B1553_FSM_Wait_RDY : constant is 1;
    attribute mti_svvh_generic_type of B1553_FSM_Over : constant is 1;
    attribute mti_svvh_generic_type of B1553_DATA_DIR_IN : constant is 1;
    attribute mti_svvh_generic_type of B1553_DATA_DIR_OUT : constant is 1;
end AHBLite_1553_Bridge;
