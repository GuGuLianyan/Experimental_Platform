library verilog;
use verilog.vl_types.all;
entity Bridge_CAN_tb is
end Bridge_CAN_tb;
