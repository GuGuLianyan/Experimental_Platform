//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Wed Mar 17 13:31:33 2021
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// SRAM_12x16
module SRAM_12x16(
    // Inputs
    CLK,
    RADDR,
    WADDR,
    WD,
    WEN,
    // Outputs
    RD
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input         CLK;
input  [3:0]  RADDR;
input  [3:0]  WADDR;
input  [11:0] WD;
input         WEN;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [11:0] RD;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire          CLK;
wire   [3:0]  RADDR;
wire   [11:0] RD_0;
wire   [3:0]  WADDR;
wire   [11:0] WD;
wire          WEN;
wire   [11:0] RD_0_net_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire          GND_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net = 1'b0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign RD_0_net_0 = RD_0;
assign RD[11:0]   = RD_0_net_0;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------SRAM_12x16_SRAM_12x16_0_TPSRAM   -   Actel:SgCore:TPSRAM:1.0.101
SRAM_12x16_SRAM_12x16_0_TPSRAM SRAM_12x16_0(
        // Inputs
        .WD    ( WD ),
        .WADDR ( WADDR ),
        .RADDR ( RADDR ),
        .WEN   ( WEN ),
        .CLK   ( CLK ),
        // Outputs
        .RD    ( RD_0 ) 
        );


endmodule
